// Emulation Verification Engineering - verilog generator
// ------------------------------------------------------
// Netlist : alb_mss_mem_lat_0000_ZMEM_i_rdel_mem   -   root module : z_alb_mss_mem_lat_0000_ZMEM_i_rdel_mem

`timescale 100 ps / 10 ps

// library : znetgen --------------------------------------------

module zview (
   I
  );
input   I;



endmodule


// library : work --------------------------------------------

module ZXLSYS (
   CLK_200
  ,CLK_100
  ,CLK_50
  ,CLK_25
  );
output  CLK_200;
output  CLK_100;
output  CLK_50;
output  CLK_25;



endmodule

module z_alb_mss_mem_lat_0000_ZMEM_i_rdel_mem (
   W0WE
  ,W0CLK
  ,W0DI
  ,W0ADDR
  ,R1DO
  ,R1ADDR
  );
input   W0WE;
input   W0CLK;
input  [130:0] W0DI;
input  [9:0] W0ADDR;
output [130:0] R1DO;
input  [9:0] R1ADDR;

wire RAMB36E1_DOBDO_0_;
wire alb_mss_mem_lat_0000_ZMEM_i_rdel_mem_add_gnd;
wire alb_mss_mem_lat_0000_ZMEM_i_rdel_mem_add_vcc;
wire RAMB36E1_0_DOBDO_0_;
wire RAMB36E1_1_DOBDO_0_;
wire RAMB36E1_2_DOBDO_0_;
wire PROTECTED_SETUP_r1addr_0_;
wire wire_sysFreq;
wire PROTECTED_SETUP_r1addr_1_;
wire PROTECTED_SETUP_r1addr_2_;
wire PROTECTED_SETUP_r1addr_3_;
wire PROTECTED_SETUP_r1addr_4_;
wire PROTECTED_SETUP_r1addr_5_;
wire PROTECTED_SETUP_r1addr_6_;
wire PROTECTED_SETUP_r1addr_7_;
wire PROTECTED_SETUP_r1addr_8_;
wire PROTECTED_SETUP_r1addr_9_;
wire w0di_0_;
wire w0di_1_;
wire w0di_2_;
wire w0di_3_;
wire w0di_4_;
wire w0di_5_;
wire w0di_6_;
wire w0di_7_;
wire w0di_8_;
wire w0di_9_;
wire w0di_10_;
wire w0di_11_;
wire w0di_12_;
wire w0di_13_;
wire w0di_14_;
wire w0di_15_;
wire w0di_16_;
wire w0di_17_;
wire w0di_18_;
wire w0di_19_;
wire w0di_20_;
wire w0di_21_;
wire w0di_22_;
wire w0di_23_;
wire w0di_24_;
wire w0di_25_;
wire w0di_26_;
wire w0di_27_;
wire w0di_28_;
wire w0di_29_;
wire w0di_30_;
wire w0di_31_;
wire w0di_32_;
wire w0di_33_;
wire w0di_34_;
wire w0di_35_;
wire w0di_36_;
wire w0di_37_;
wire w0di_38_;
wire w0di_39_;
wire w0di_40_;
wire w0di_41_;
wire w0di_42_;
wire w0di_43_;
wire w0di_44_;
wire w0di_45_;
wire w0di_46_;
wire w0di_47_;
wire w0di_48_;
wire w0di_49_;
wire w0di_50_;
wire w0di_51_;
wire w0di_52_;
wire w0di_53_;
wire w0di_54_;
wire w0di_55_;
wire w0di_56_;
wire w0di_57_;
wire w0di_58_;
wire w0di_59_;
wire w0di_60_;
wire w0di_61_;
wire w0di_62_;
wire w0di_63_;
wire w0di_64_;
wire w0di_65_;
wire w0di_66_;
wire w0di_67_;
wire w0di_68_;
wire w0di_69_;
wire w0di_70_;
wire w0di_71_;
wire w0di_72_;
wire w0di_73_;
wire w0di_74_;
wire w0di_75_;
wire w0di_76_;
wire w0di_77_;
wire w0di_78_;
wire w0di_79_;
wire w0di_80_;
wire w0di_81_;
wire w0di_82_;
wire w0di_83_;
wire w0di_84_;
wire w0di_85_;
wire w0di_86_;
wire w0di_87_;
wire w0di_88_;
wire w0di_89_;
wire w0di_90_;
wire w0di_91_;
wire w0di_92_;
wire w0di_93_;
wire w0di_94_;
wire w0di_95_;
wire w0di_96_;
wire w0di_97_;
wire w0di_98_;
wire w0di_99_;
wire w0di_100_;
wire w0di_101_;
wire w0di_102_;
wire w0di_103_;
wire w0di_104_;
wire w0di_105_;
wire w0di_106_;
wire w0di_107_;
wire w0di_108_;
wire w0di_109_;
wire w0di_110_;
wire w0di_111_;
wire w0di_112_;
wire w0di_113_;
wire w0di_114_;
wire w0di_115_;
wire w0di_116_;
wire w0di_117_;
wire w0di_118_;
wire w0di_119_;
wire w0di_120_;
wire w0di_121_;
wire w0di_122_;
wire w0di_123_;
wire w0di_124_;
wire w0di_125_;
wire w0di_126_;
wire w0di_127_;
wire w0di_128_;
wire w0di_129_;
wire w0di_130_;
wire w0we;
wire w0clk;
wire w0addr_0_;
wire w0addr_1_;
wire w0addr_2_;
wire w0addr_3_;
wire w0addr_4_;
wire w0addr_5_;
wire w0addr_6_;
wire w0addr_7_;
wire w0addr_8_;
wire w0addr_9_;
wire r1do_0_;
wire r1do_1_;
wire r1do_2_;
wire r1do_3_;
wire r1do_4_;
wire r1do_5_;
wire r1do_6_;
wire r1do_7_;
wire r1do_8_;
wire r1do_9_;
wire r1do_10_;
wire r1do_11_;
wire r1do_12_;
wire r1do_13_;
wire r1do_14_;
wire r1do_15_;
wire r1do_16_;
wire r1do_17_;
wire r1do_18_;
wire r1do_19_;
wire r1do_20_;
wire r1do_21_;
wire r1do_22_;
wire r1do_23_;
wire r1do_24_;
wire r1do_25_;
wire r1do_26_;
wire r1do_27_;
wire r1do_28_;
wire r1do_29_;
wire r1do_30_;
wire r1do_31_;
wire r1do_32_;
wire r1do_33_;
wire r1do_34_;
wire r1do_35_;
wire r1do_36_;
wire r1do_37_;
wire r1do_38_;
wire r1do_39_;
wire r1do_40_;
wire r1do_41_;
wire r1do_42_;
wire r1do_43_;
wire r1do_44_;
wire r1do_45_;
wire r1do_46_;
wire r1do_47_;
wire r1do_48_;
wire r1do_49_;
wire r1do_50_;
wire r1do_51_;
wire r1do_52_;
wire r1do_53_;
wire r1do_54_;
wire r1do_55_;
wire r1do_56_;
wire r1do_57_;
wire r1do_58_;
wire r1do_59_;
wire r1do_60_;
wire r1do_61_;
wire r1do_62_;
wire r1do_63_;
wire r1do_64_;
wire r1do_65_;
wire r1do_66_;
wire r1do_67_;
wire r1do_68_;
wire r1do_69_;
wire r1do_70_;
wire r1do_71_;
wire r1do_72_;
wire r1do_73_;
wire r1do_74_;
wire r1do_75_;
wire r1do_76_;
wire r1do_77_;
wire r1do_78_;
wire r1do_79_;
wire r1do_80_;
wire r1do_81_;
wire r1do_82_;
wire r1do_83_;
wire r1do_84_;
wire r1do_85_;
wire r1do_86_;
wire r1do_87_;
wire r1do_88_;
wire r1do_89_;
wire r1do_90_;
wire r1do_91_;
wire r1do_92_;
wire r1do_93_;
wire r1do_94_;
wire r1do_95_;
wire r1do_96_;
wire r1do_97_;
wire r1do_98_;
wire r1do_99_;
wire r1do_100_;
wire r1do_101_;
wire r1do_102_;
wire r1do_103_;
wire r1do_104_;
wire r1do_105_;
wire r1do_106_;
wire r1do_107_;
wire r1do_108_;
wire r1do_109_;
wire r1do_110_;
wire r1do_111_;
wire r1do_112_;
wire r1do_113_;
wire r1do_114_;
wire r1do_115_;
wire r1do_116_;
wire r1do_117_;
wire r1do_118_;
wire r1do_119_;
wire r1do_120_;
wire r1do_121_;
wire r1do_122_;
wire r1do_123_;
wire r1do_124_;
wire r1do_125_;
wire r1do_126_;
wire r1do_127_;
wire r1do_128_;
wire r1do_129_;
wire r1do_130_;
wire r1addr_0_;
wire r1addr_1_;
wire r1addr_2_;
wire r1addr_3_;
wire r1addr_4_;
wire r1addr_5_;
wire r1addr_6_;
wire r1addr_7_;
wire r1addr_8_;
wire r1addr_9_;
wire zsimv_ucon_0;
wire zsimv_ucon_1;
wire zsimv_ucon_2;
wire zsimv_ucon_3;
wire zsimv_ucon_4;
wire zsimv_ucon_5;
wire zsimv_ucon_6;
wire zsimv_ucon_7;
wire zsimv_ucon_8;
wire zsimv_ucon_9;
wire zsimv_ucon_10;
wire zsimv_ucon_11;
wire zsimv_ucon_12;
wire zsimv_ucon_13;
wire zsimv_ucon_14;
wire zsimv_ucon_15;
wire zsimv_ucon_16;
wire zsimv_ucon_17;
wire zsimv_ucon_18;
wire zsimv_ucon_19;
wire zsimv_ucon_20;
wire zsimv_ucon_21;
wire zsimv_ucon_22;
wire zsimv_ucon_23;
wire zsimv_ucon_24;
wire zsimv_ucon_25;
wire zsimv_ucon_26;
wire zsimv_ucon_27;
wire zsimv_ucon_28;
wire zsimv_ucon_29;
wire zsimv_ucon_30;
wire zsimv_ucon_31;
wire zsimv_ucon_32;
wire zsimv_ucon_33;
wire zsimv_ucon_34;
wire zsimv_ucon_35;
wire zsimv_ucon_36;
wire zsimv_ucon_37;
wire zsimv_ucon_38;
wire zsimv_ucon_39;
wire zsimv_ucon_40;
wire zsimv_ucon_41;
wire zsimv_ucon_42;
wire zsimv_ucon_43;
wire zsimv_ucon_44;
wire zsimv_ucon_45;
wire zsimv_ucon_46;
wire zsimv_ucon_47;
wire zsimv_ucon_48;
wire zsimv_ucon_49;
wire zsimv_ucon_50;
wire zsimv_ucon_51;
wire zsimv_ucon_52;
wire zsimv_ucon_53;
wire zsimv_ucon_54;
wire zsimv_ucon_55;
wire zsimv_ucon_56;
wire zsimv_ucon_57;
wire zsimv_ucon_58;
wire zsimv_ucon_59;
wire zsimv_ucon_60;
wire zsimv_ucon_61;
wire zsimv_ucon_62;
wire zsimv_ucon_63;
wire zsimv_ucon_64;
wire zsimv_ucon_65;
wire zsimv_ucon_66;
wire zsimv_ucon_67;
wire zsimv_ucon_68;
wire zsimv_ucon_69;
wire zsimv_ucon_70;
wire zsimv_ucon_71;
wire zsimv_ucon_72;
wire zsimv_ucon_73;
wire zsimv_ucon_74;
wire zsimv_ucon_75;
wire zsimv_ucon_76;
wire zsimv_ucon_77;
wire zsimv_ucon_78;
wire zsimv_ucon_79;
wire zsimv_ucon_80;
wire zsimv_ucon_81;
wire zsimv_ucon_82;
wire zsimv_ucon_83;
wire zsimv_ucon_84;
wire zsimv_ucon_85;
wire zsimv_ucon_86;
wire zsimv_ucon_87;
wire zsimv_ucon_88;
wire zsimv_ucon_89;
wire zsimv_ucon_90;
wire zsimv_ucon_91;
wire zsimv_ucon_92;
wire zsimv_ucon_93;
wire zsimv_ucon_94;
wire zsimv_ucon_95;
wire zsimv_ucon_96;
wire zsimv_ucon_97;
wire zsimv_ucon_98;
wire zsimv_ucon_99;
wire zsimv_ucon_100;
wire zsimv_ucon_101;
wire zsimv_ucon_102;
wire zsimv_ucon_103;
wire zsimv_ucon_104;
wire zsimv_ucon_105;
wire zsimv_ucon_106;
wire zsimv_ucon_107;
wire zsimv_ucon_108;
wire zsimv_ucon_109;
wire zsimv_ucon_110;
wire zsimv_ucon_111;
wire zsimv_ucon_112;
wire zsimv_ucon_113;
wire zsimv_ucon_114;
wire zsimv_ucon_115;
wire zsimv_ucon_116;
wire zsimv_ucon_117;
wire zsimv_ucon_118;
wire zsimv_ucon_119;
wire zsimv_ucon_120;
wire zsimv_ucon_121;
wire zsimv_ucon_122;
wire zsimv_ucon_123;
wire zsimv_ucon_124;
wire zsimv_ucon_125;
wire zsimv_ucon_126;
wire zsimv_ucon_127;
wire zsimv_ucon_128;
wire zsimv_ucon_129;
wire zsimv_ucon_130;
wire zsimv_ucon_131;
wire zsimv_ucon_132;
wire zsimv_ucon_133;
wire zsimv_ucon_134;
wire zsimv_ucon_135;
wire zsimv_ucon_136;
wire zsimv_ucon_137;
wire zsimv_ucon_138;
wire zsimv_ucon_139;
wire zsimv_ucon_140;
wire zsimv_ucon_141;
wire zsimv_ucon_142;
wire zsimv_ucon_143;
wire zsimv_ucon_144;
wire zsimv_ucon_145;
wire zsimv_ucon_146;
wire zsimv_ucon_147;
wire zsimv_ucon_148;
wire zsimv_ucon_149;
wire zsimv_ucon_150;
wire zsimv_ucon_151;
wire zsimv_ucon_152;
wire zsimv_ucon_153;
wire zsimv_ucon_154;
wire zsimv_ucon_155;
wire zsimv_ucon_156;
wire zsimv_ucon_157;
wire zsimv_ucon_158;
wire zsimv_ucon_159;
wire zsimv_ucon_160;
wire zsimv_ucon_161;
wire zsimv_ucon_162;
wire zsimv_ucon_163;
wire zsimv_ucon_164;
wire zsimv_ucon_165;
wire zsimv_ucon_166;
wire zsimv_ucon_167;
wire zsimv_ucon_168;
wire zsimv_ucon_169;
wire zsimv_ucon_170;
wire zsimv_ucon_171;
wire zsimv_ucon_172;
wire zsimv_ucon_173;
wire zsimv_ucon_174;
wire zsimv_ucon_175;
wire zsimv_ucon_176;
wire zsimv_ucon_177;
wire zsimv_ucon_178;
wire zsimv_ucon_179;
wire zsimv_ucon_180;
wire zsimv_ucon_181;
wire zsimv_ucon_182;
wire zsimv_ucon_183;
wire zsimv_ucon_184;
wire zsimv_ucon_185;
wire zsimv_ucon_186;
wire zsimv_ucon_187;
wire zsimv_ucon_188;
wire zsimv_ucon_189;
wire zsimv_ucon_190;
wire zsimv_ucon_191;
wire zsimv_ucon_192;
wire zsimv_ucon_193;
wire zsimv_ucon_194;
wire zsimv_ucon_195;
wire zsimv_ucon_196;
wire zsimv_ucon_197;
wire zsimv_ucon_198;
wire zsimv_ucon_199;
wire zsimv_ucon_200;
wire zsimv_ucon_201;
wire zsimv_ucon_202;
wire zsimv_ucon_203;
wire zsimv_ucon_204;
wire zsimv_ucon_205;
wire zsimv_ucon_206;
wire zsimv_ucon_207;
wire zsimv_ucon_208;
wire zsimv_ucon_209;
wire zsimv_ucon_210;
wire zsimv_ucon_211;
wire zsimv_ucon_212;
wire zsimv_ucon_213;
wire zsimv_ucon_214;
wire zsimv_ucon_215;
wire zsimv_ucon_216;
wire zsimv_ucon_217;
wire zsimv_ucon_218;
wire zsimv_ucon_219;
wire zsimv_ucon_220;
wire zsimv_ucon_221;
wire zsimv_ucon_222;
wire zsimv_ucon_223;
wire zsimv_ucon_224;
wire zsimv_ucon_225;
wire zsimv_ucon_226;
wire zsimv_ucon_227;
wire zsimv_ucon_228;
wire zsimv_ucon_229;
wire zsimv_ucon_230;
wire zsimv_ucon_231;
wire zsimv_ucon_232;
wire zsimv_ucon_233;
wire zsimv_ucon_234;
wire zsimv_ucon_235;
wire zsimv_ucon_236;
wire zsimv_ucon_237;
wire zsimv_ucon_238;
wire zsimv_ucon_239;
wire zsimv_ucon_240;
wire zsimv_ucon_241;
wire zsimv_ucon_242;
wire zsimv_ucon_243;
wire zsimv_ucon_244;
wire zsimv_ucon_245;
wire zsimv_ucon_246;
wire zsimv_ucon_247;
wire zsimv_ucon_248;
wire zsimv_ucon_249;
wire zsimv_ucon_250;
wire zsimv_ucon_251;
wire zsimv_ucon_252;
wire zsimv_ucon_253;
wire zsimv_ucon_254;
wire zsimv_ucon_255;

assign w0di_0_ = W0DI[0];
assign w0di_1_ = W0DI[1];
assign w0di_2_ = W0DI[2];
assign w0di_3_ = W0DI[3];
assign w0di_4_ = W0DI[4];
assign w0di_5_ = W0DI[5];
assign w0di_6_ = W0DI[6];
assign w0di_7_ = W0DI[7];
assign w0di_8_ = W0DI[8];
assign w0di_9_ = W0DI[9];
assign w0di_10_ = W0DI[10];
assign w0di_11_ = W0DI[11];
assign w0di_12_ = W0DI[12];
assign w0di_13_ = W0DI[13];
assign w0di_14_ = W0DI[14];
assign w0di_15_ = W0DI[15];
assign w0di_16_ = W0DI[16];
assign w0di_17_ = W0DI[17];
assign w0di_18_ = W0DI[18];
assign w0di_19_ = W0DI[19];
assign w0di_20_ = W0DI[20];
assign w0di_21_ = W0DI[21];
assign w0di_22_ = W0DI[22];
assign w0di_23_ = W0DI[23];
assign w0di_24_ = W0DI[24];
assign w0di_25_ = W0DI[25];
assign w0di_26_ = W0DI[26];
assign w0di_27_ = W0DI[27];
assign w0di_28_ = W0DI[28];
assign w0di_29_ = W0DI[29];
assign w0di_30_ = W0DI[30];
assign w0di_31_ = W0DI[31];
assign w0di_32_ = W0DI[32];
assign w0di_33_ = W0DI[33];
assign w0di_34_ = W0DI[34];
assign w0di_35_ = W0DI[35];
assign w0di_36_ = W0DI[36];
assign w0di_37_ = W0DI[37];
assign w0di_38_ = W0DI[38];
assign w0di_39_ = W0DI[39];
assign w0di_40_ = W0DI[40];
assign w0di_41_ = W0DI[41];
assign w0di_42_ = W0DI[42];
assign w0di_43_ = W0DI[43];
assign w0di_44_ = W0DI[44];
assign w0di_45_ = W0DI[45];
assign w0di_46_ = W0DI[46];
assign w0di_47_ = W0DI[47];
assign w0di_48_ = W0DI[48];
assign w0di_49_ = W0DI[49];
assign w0di_50_ = W0DI[50];
assign w0di_51_ = W0DI[51];
assign w0di_52_ = W0DI[52];
assign w0di_53_ = W0DI[53];
assign w0di_54_ = W0DI[54];
assign w0di_55_ = W0DI[55];
assign w0di_56_ = W0DI[56];
assign w0di_57_ = W0DI[57];
assign w0di_58_ = W0DI[58];
assign w0di_59_ = W0DI[59];
assign w0di_60_ = W0DI[60];
assign w0di_61_ = W0DI[61];
assign w0di_62_ = W0DI[62];
assign w0di_63_ = W0DI[63];
assign w0di_64_ = W0DI[64];
assign w0di_65_ = W0DI[65];
assign w0di_66_ = W0DI[66];
assign w0di_67_ = W0DI[67];
assign w0di_68_ = W0DI[68];
assign w0di_69_ = W0DI[69];
assign w0di_70_ = W0DI[70];
assign w0di_71_ = W0DI[71];
assign w0di_72_ = W0DI[72];
assign w0di_73_ = W0DI[73];
assign w0di_74_ = W0DI[74];
assign w0di_75_ = W0DI[75];
assign w0di_76_ = W0DI[76];
assign w0di_77_ = W0DI[77];
assign w0di_78_ = W0DI[78];
assign w0di_79_ = W0DI[79];
assign w0di_80_ = W0DI[80];
assign w0di_81_ = W0DI[81];
assign w0di_82_ = W0DI[82];
assign w0di_83_ = W0DI[83];
assign w0di_84_ = W0DI[84];
assign w0di_85_ = W0DI[85];
assign w0di_86_ = W0DI[86];
assign w0di_87_ = W0DI[87];
assign w0di_88_ = W0DI[88];
assign w0di_89_ = W0DI[89];
assign w0di_90_ = W0DI[90];
assign w0di_91_ = W0DI[91];
assign w0di_92_ = W0DI[92];
assign w0di_93_ = W0DI[93];
assign w0di_94_ = W0DI[94];
assign w0di_95_ = W0DI[95];
assign w0di_96_ = W0DI[96];
assign w0di_97_ = W0DI[97];
assign w0di_98_ = W0DI[98];
assign w0di_99_ = W0DI[99];
assign w0di_100_ = W0DI[100];
assign w0di_101_ = W0DI[101];
assign w0di_102_ = W0DI[102];
assign w0di_103_ = W0DI[103];
assign w0di_104_ = W0DI[104];
assign w0di_105_ = W0DI[105];
assign w0di_106_ = W0DI[106];
assign w0di_107_ = W0DI[107];
assign w0di_108_ = W0DI[108];
assign w0di_109_ = W0DI[109];
assign w0di_110_ = W0DI[110];
assign w0di_111_ = W0DI[111];
assign w0di_112_ = W0DI[112];
assign w0di_113_ = W0DI[113];
assign w0di_114_ = W0DI[114];
assign w0di_115_ = W0DI[115];
assign w0di_116_ = W0DI[116];
assign w0di_117_ = W0DI[117];
assign w0di_118_ = W0DI[118];
assign w0di_119_ = W0DI[119];
assign w0di_120_ = W0DI[120];
assign w0di_121_ = W0DI[121];
assign w0di_122_ = W0DI[122];
assign w0di_123_ = W0DI[123];
assign w0di_124_ = W0DI[124];
assign w0di_125_ = W0DI[125];
assign w0di_126_ = W0DI[126];
assign w0di_127_ = W0DI[127];
assign w0di_128_ = W0DI[128];
assign w0di_129_ = W0DI[129];
assign w0di_130_ = W0DI[130];
assign w0we = W0WE;
assign w0clk = W0CLK;
assign w0addr_0_ = W0ADDR[0];
assign w0addr_1_ = W0ADDR[1];
assign w0addr_2_ = W0ADDR[2];
assign w0addr_3_ = W0ADDR[3];
assign w0addr_4_ = W0ADDR[4];
assign w0addr_5_ = W0ADDR[5];
assign w0addr_6_ = W0ADDR[6];
assign w0addr_7_ = W0ADDR[7];
assign w0addr_8_ = W0ADDR[8];
assign w0addr_9_ = W0ADDR[9];
assign R1DO[0] = r1do_0_;
assign R1DO[1] = r1do_1_;
assign R1DO[2] = r1do_2_;
assign R1DO[3] = r1do_3_;
assign R1DO[4] = r1do_4_;
assign R1DO[5] = r1do_5_;
assign R1DO[6] = r1do_6_;
assign R1DO[7] = r1do_7_;
assign R1DO[8] = r1do_8_;
assign R1DO[9] = r1do_9_;
assign R1DO[10] = r1do_10_;
assign R1DO[11] = r1do_11_;
assign R1DO[12] = r1do_12_;
assign R1DO[13] = r1do_13_;
assign R1DO[14] = r1do_14_;
assign R1DO[15] = r1do_15_;
assign R1DO[16] = r1do_16_;
assign R1DO[17] = r1do_17_;
assign R1DO[18] = r1do_18_;
assign R1DO[19] = r1do_19_;
assign R1DO[20] = r1do_20_;
assign R1DO[21] = r1do_21_;
assign R1DO[22] = r1do_22_;
assign R1DO[23] = r1do_23_;
assign R1DO[24] = r1do_24_;
assign R1DO[25] = r1do_25_;
assign R1DO[26] = r1do_26_;
assign R1DO[27] = r1do_27_;
assign R1DO[28] = r1do_28_;
assign R1DO[29] = r1do_29_;
assign R1DO[30] = r1do_30_;
assign R1DO[31] = r1do_31_;
assign R1DO[32] = r1do_32_;
assign R1DO[33] = r1do_33_;
assign R1DO[34] = r1do_34_;
assign R1DO[35] = r1do_35_;
assign R1DO[36] = r1do_36_;
assign R1DO[37] = r1do_37_;
assign R1DO[38] = r1do_38_;
assign R1DO[39] = r1do_39_;
assign R1DO[40] = r1do_40_;
assign R1DO[41] = r1do_41_;
assign R1DO[42] = r1do_42_;
assign R1DO[43] = r1do_43_;
assign R1DO[44] = r1do_44_;
assign R1DO[45] = r1do_45_;
assign R1DO[46] = r1do_46_;
assign R1DO[47] = r1do_47_;
assign R1DO[48] = r1do_48_;
assign R1DO[49] = r1do_49_;
assign R1DO[50] = r1do_50_;
assign R1DO[51] = r1do_51_;
assign R1DO[52] = r1do_52_;
assign R1DO[53] = r1do_53_;
assign R1DO[54] = r1do_54_;
assign R1DO[55] = r1do_55_;
assign R1DO[56] = r1do_56_;
assign R1DO[57] = r1do_57_;
assign R1DO[58] = r1do_58_;
assign R1DO[59] = r1do_59_;
assign R1DO[60] = r1do_60_;
assign R1DO[61] = r1do_61_;
assign R1DO[62] = r1do_62_;
assign R1DO[63] = r1do_63_;
assign R1DO[64] = r1do_64_;
assign R1DO[65] = r1do_65_;
assign R1DO[66] = r1do_66_;
assign R1DO[67] = r1do_67_;
assign R1DO[68] = r1do_68_;
assign R1DO[69] = r1do_69_;
assign R1DO[70] = r1do_70_;
assign R1DO[71] = r1do_71_;
assign R1DO[72] = r1do_72_;
assign R1DO[73] = r1do_73_;
assign R1DO[74] = r1do_74_;
assign R1DO[75] = r1do_75_;
assign R1DO[76] = r1do_76_;
assign R1DO[77] = r1do_77_;
assign R1DO[78] = r1do_78_;
assign R1DO[79] = r1do_79_;
assign R1DO[80] = r1do_80_;
assign R1DO[81] = r1do_81_;
assign R1DO[82] = r1do_82_;
assign R1DO[83] = r1do_83_;
assign R1DO[84] = r1do_84_;
assign R1DO[85] = r1do_85_;
assign R1DO[86] = r1do_86_;
assign R1DO[87] = r1do_87_;
assign R1DO[88] = r1do_88_;
assign R1DO[89] = r1do_89_;
assign R1DO[90] = r1do_90_;
assign R1DO[91] = r1do_91_;
assign R1DO[92] = r1do_92_;
assign R1DO[93] = r1do_93_;
assign R1DO[94] = r1do_94_;
assign R1DO[95] = r1do_95_;
assign R1DO[96] = r1do_96_;
assign R1DO[97] = r1do_97_;
assign R1DO[98] = r1do_98_;
assign R1DO[99] = r1do_99_;
assign R1DO[100] = r1do_100_;
assign R1DO[101] = r1do_101_;
assign R1DO[102] = r1do_102_;
assign R1DO[103] = r1do_103_;
assign R1DO[104] = r1do_104_;
assign R1DO[105] = r1do_105_;
assign R1DO[106] = r1do_106_;
assign R1DO[107] = r1do_107_;
assign R1DO[108] = r1do_108_;
assign R1DO[109] = r1do_109_;
assign R1DO[110] = r1do_110_;
assign R1DO[111] = r1do_111_;
assign R1DO[112] = r1do_112_;
assign R1DO[113] = r1do_113_;
assign R1DO[114] = r1do_114_;
assign R1DO[115] = r1do_115_;
assign R1DO[116] = r1do_116_;
assign R1DO[117] = r1do_117_;
assign R1DO[118] = r1do_118_;
assign R1DO[119] = r1do_119_;
assign R1DO[120] = r1do_120_;
assign R1DO[121] = r1do_121_;
assign R1DO[122] = r1do_122_;
assign R1DO[123] = r1do_123_;
assign R1DO[124] = r1do_124_;
assign R1DO[125] = r1do_125_;
assign R1DO[126] = r1do_126_;
assign R1DO[127] = r1do_127_;
assign R1DO[128] = r1do_128_;
assign R1DO[129] = r1do_129_;
assign R1DO[130] = r1do_130_;
assign r1addr_0_ = R1ADDR[0];
assign r1addr_1_ = R1ADDR[1];
assign r1addr_2_ = R1ADDR[2];
assign r1addr_3_ = R1ADDR[3];
assign r1addr_4_ = R1ADDR[4];
assign r1addr_5_ = R1ADDR[5];
assign r1addr_6_ = R1ADDR[6];
assign r1addr_7_ = R1ADDR[7];
assign r1addr_8_ = R1ADDR[8];
assign r1addr_9_ = R1ADDR[9];

GND I_alb_mss_mem_lat_0000_ZMEM_i_rdel_mem_add_gnd (
    .G(alb_mss_mem_lat_0000_ZMEM_i_rdel_mem_add_gnd)
  );

VCC I_alb_mss_mem_lat_0000_ZMEM_i_rdel_mem_add_vcc (
    .P(alb_mss_mem_lat_0000_ZMEM_i_rdel_mem_add_vcc)
  );

FD \I_PROTECTED_SETUP_r1addr[0]  (
    .Q(PROTECTED_SETUP_r1addr_0_)
  , .C(wire_sysFreq)
  , .D(r1addr_0_)
  );

ZXLSYS I_zgatezxlsys (
    .CLK_200(zsimv_ucon_0)
  , .CLK_100(wire_sysFreq)
  , .CLK_50(zsimv_ucon_1)
  , .CLK_25(zsimv_ucon_2)
  );

FD \I_PROTECTED_SETUP_r1addr[1]  (
    .Q(PROTECTED_SETUP_r1addr_1_)
  , .C(wire_sysFreq)
  , .D(r1addr_1_)
  );

FD \I_PROTECTED_SETUP_r1addr[2]  (
    .Q(PROTECTED_SETUP_r1addr_2_)
  , .C(wire_sysFreq)
  , .D(r1addr_2_)
  );

FD \I_PROTECTED_SETUP_r1addr[3]  (
    .Q(PROTECTED_SETUP_r1addr_3_)
  , .C(wire_sysFreq)
  , .D(r1addr_3_)
  );

FD \I_PROTECTED_SETUP_r1addr[4]  (
    .Q(PROTECTED_SETUP_r1addr_4_)
  , .C(wire_sysFreq)
  , .D(r1addr_4_)
  );

FD \I_PROTECTED_SETUP_r1addr[5]  (
    .Q(PROTECTED_SETUP_r1addr_5_)
  , .C(wire_sysFreq)
  , .D(r1addr_5_)
  );

FD \I_PROTECTED_SETUP_r1addr[6]  (
    .Q(PROTECTED_SETUP_r1addr_6_)
  , .C(wire_sysFreq)
  , .D(r1addr_6_)
  );

FD \I_PROTECTED_SETUP_r1addr[7]  (
    .Q(PROTECTED_SETUP_r1addr_7_)
  , .C(wire_sysFreq)
  , .D(r1addr_7_)
  );

FD \I_PROTECTED_SETUP_r1addr[8]  (
    .Q(PROTECTED_SETUP_r1addr_8_)
  , .C(wire_sysFreq)
  , .D(r1addr_8_)
  );

FD \I_PROTECTED_SETUP_r1addr[9]  (
    .Q(PROTECTED_SETUP_r1addr_9_)
  , .C(wire_sysFreq)
  , .D(r1addr_9_)
  );

defparam I_RAMB36E1.SRVAL_A = "000000000000000000000000000000000000";
defparam I_RAMB36E1.SRVAL_B = "000000000000000000000000000000000000";
defparam I_RAMB36E1.WRITE_MODE_A = "READ_FIRST";
defparam I_RAMB36E1.WRITE_MODE_B = "READ_FIRST";
defparam I_RAMB36E1.WRITE_WIDTH_B = 36;
defparam I_RAMB36E1.READ_WIDTH_A = 36;
RAMB36E1 I_RAMB36E1 (
    .CASCADEOUTA(zsimv_ucon_3)
  , .CASCADEOUTB(zsimv_ucon_4)
  , .DBITERR(zsimv_ucon_5)
  , .SBITERR(zsimv_ucon_58)
  , .CASCADEINA(zsimv_ucon_59)
  , .CASCADEINB(zsimv_ucon_60)
  , .CLKARDCLK(wire_sysFreq)
  , .CLKBWRCLK(w0clk)
  , .ENARDEN(alb_mss_mem_lat_0000_ZMEM_i_rdel_mem_add_vcc)
  , .ENBWREN(alb_mss_mem_lat_0000_ZMEM_i_rdel_mem_add_vcc)
  , .INJECTDBITERR(zsimv_ucon_61)
  , .INJECTSBITERR(zsimv_ucon_62)
  , .REGCEAREGCE(alb_mss_mem_lat_0000_ZMEM_i_rdel_mem_add_gnd)
  , .REGCEB(alb_mss_mem_lat_0000_ZMEM_i_rdel_mem_add_gnd)
  , .RSTRAMARSTRAM(alb_mss_mem_lat_0000_ZMEM_i_rdel_mem_add_gnd)
  , .RSTRAMB(alb_mss_mem_lat_0000_ZMEM_i_rdel_mem_add_gnd)
  , .RSTREGARSTREG(alb_mss_mem_lat_0000_ZMEM_i_rdel_mem_add_gnd)
  , .RSTREGB(alb_mss_mem_lat_0000_ZMEM_i_rdel_mem_add_gnd)
  , .DIPADIP(
   {  alb_mss_mem_lat_0000_ZMEM_i_rdel_mem_add_gnd, alb_mss_mem_lat_0000_ZMEM_i_rdel_mem_add_gnd, alb_mss_mem_lat_0000_ZMEM_i_rdel_mem_add_gnd, alb_mss_mem_lat_0000_ZMEM_i_rdel_mem_add_gnd
   } )
  , .DIPBDIP(
   {  w0di_35_, w0di_34_, w0di_33_, w0di_32_
   } )
  , .WEA(
   {  alb_mss_mem_lat_0000_ZMEM_i_rdel_mem_add_gnd, alb_mss_mem_lat_0000_ZMEM_i_rdel_mem_add_gnd, alb_mss_mem_lat_0000_ZMEM_i_rdel_mem_add_gnd, alb_mss_mem_lat_0000_ZMEM_i_rdel_mem_add_gnd
   } )
  , .WEBWE(
   {  w0we, w0we, w0we, w0we
  , w0we, w0we, w0we, w0we
   } )
  , .ADDRARDADDR(
   {  alb_mss_mem_lat_0000_ZMEM_i_rdel_mem_add_gnd, PROTECTED_SETUP_r1addr_9_, PROTECTED_SETUP_r1addr_8_, PROTECTED_SETUP_r1addr_7_
  , PROTECTED_SETUP_r1addr_6_, PROTECTED_SETUP_r1addr_5_, PROTECTED_SETUP_r1addr_4_, PROTECTED_SETUP_r1addr_3_
  , PROTECTED_SETUP_r1addr_2_, PROTECTED_SETUP_r1addr_1_, PROTECTED_SETUP_r1addr_0_, alb_mss_mem_lat_0000_ZMEM_i_rdel_mem_add_gnd
  , alb_mss_mem_lat_0000_ZMEM_i_rdel_mem_add_gnd, alb_mss_mem_lat_0000_ZMEM_i_rdel_mem_add_gnd, alb_mss_mem_lat_0000_ZMEM_i_rdel_mem_add_gnd, alb_mss_mem_lat_0000_ZMEM_i_rdel_mem_add_gnd
   } )
  , .ADDRBWRADDR(
   {  alb_mss_mem_lat_0000_ZMEM_i_rdel_mem_add_gnd, w0addr_9_, w0addr_8_, w0addr_7_
  , w0addr_6_, w0addr_5_, w0addr_4_, w0addr_3_
  , w0addr_2_, w0addr_1_, w0addr_0_, alb_mss_mem_lat_0000_ZMEM_i_rdel_mem_add_gnd
  , alb_mss_mem_lat_0000_ZMEM_i_rdel_mem_add_gnd, alb_mss_mem_lat_0000_ZMEM_i_rdel_mem_add_gnd, alb_mss_mem_lat_0000_ZMEM_i_rdel_mem_add_gnd, alb_mss_mem_lat_0000_ZMEM_i_rdel_mem_add_gnd
   } )
  , .DIADI(
   {  alb_mss_mem_lat_0000_ZMEM_i_rdel_mem_add_gnd, alb_mss_mem_lat_0000_ZMEM_i_rdel_mem_add_gnd, alb_mss_mem_lat_0000_ZMEM_i_rdel_mem_add_gnd, alb_mss_mem_lat_0000_ZMEM_i_rdel_mem_add_gnd
  , alb_mss_mem_lat_0000_ZMEM_i_rdel_mem_add_gnd, alb_mss_mem_lat_0000_ZMEM_i_rdel_mem_add_gnd, alb_mss_mem_lat_0000_ZMEM_i_rdel_mem_add_gnd, alb_mss_mem_lat_0000_ZMEM_i_rdel_mem_add_gnd
  , alb_mss_mem_lat_0000_ZMEM_i_rdel_mem_add_gnd, alb_mss_mem_lat_0000_ZMEM_i_rdel_mem_add_gnd, alb_mss_mem_lat_0000_ZMEM_i_rdel_mem_add_gnd, alb_mss_mem_lat_0000_ZMEM_i_rdel_mem_add_gnd
  , alb_mss_mem_lat_0000_ZMEM_i_rdel_mem_add_gnd, alb_mss_mem_lat_0000_ZMEM_i_rdel_mem_add_gnd, alb_mss_mem_lat_0000_ZMEM_i_rdel_mem_add_gnd, alb_mss_mem_lat_0000_ZMEM_i_rdel_mem_add_gnd
  , alb_mss_mem_lat_0000_ZMEM_i_rdel_mem_add_gnd, alb_mss_mem_lat_0000_ZMEM_i_rdel_mem_add_gnd, alb_mss_mem_lat_0000_ZMEM_i_rdel_mem_add_gnd, alb_mss_mem_lat_0000_ZMEM_i_rdel_mem_add_gnd
  , alb_mss_mem_lat_0000_ZMEM_i_rdel_mem_add_gnd, alb_mss_mem_lat_0000_ZMEM_i_rdel_mem_add_gnd, alb_mss_mem_lat_0000_ZMEM_i_rdel_mem_add_gnd, alb_mss_mem_lat_0000_ZMEM_i_rdel_mem_add_gnd
  , alb_mss_mem_lat_0000_ZMEM_i_rdel_mem_add_gnd, alb_mss_mem_lat_0000_ZMEM_i_rdel_mem_add_gnd, alb_mss_mem_lat_0000_ZMEM_i_rdel_mem_add_gnd, alb_mss_mem_lat_0000_ZMEM_i_rdel_mem_add_gnd
  , alb_mss_mem_lat_0000_ZMEM_i_rdel_mem_add_gnd, alb_mss_mem_lat_0000_ZMEM_i_rdel_mem_add_gnd, alb_mss_mem_lat_0000_ZMEM_i_rdel_mem_add_gnd, alb_mss_mem_lat_0000_ZMEM_i_rdel_mem_add_gnd
   } )
  , .DIBDI(
   {  w0di_31_, w0di_30_, w0di_29_, w0di_28_
  , w0di_27_, w0di_26_, w0di_25_, w0di_24_
  , w0di_23_, w0di_22_, w0di_21_, w0di_20_
  , w0di_19_, w0di_18_, w0di_17_, w0di_16_
  , w0di_15_, w0di_14_, w0di_13_, w0di_12_
  , w0di_11_, w0di_10_, w0di_9_, w0di_8_
  , w0di_7_, w0di_6_, w0di_5_, w0di_4_
  , w0di_3_, w0di_2_, w0di_1_, w0di_0_
   } )
  , .DOPADOP(
   {  r1do_35_, r1do_34_, r1do_33_, r1do_32_
   } )
  , .DOPBDOP(
   {  zsimv_ucon_40, zsimv_ucon_39, zsimv_ucon_38, zsimv_ucon_37
   } )
  , .ECCPARITY(
   {  zsimv_ucon_48, zsimv_ucon_47, zsimv_ucon_46, zsimv_ucon_45
  , zsimv_ucon_44, zsimv_ucon_43, zsimv_ucon_42, zsimv_ucon_41
   } )
  , .RDADDRECC(
   {  zsimv_ucon_57, zsimv_ucon_56, zsimv_ucon_55, zsimv_ucon_54
  , zsimv_ucon_53, zsimv_ucon_52, zsimv_ucon_51, zsimv_ucon_50
  , zsimv_ucon_49 } )
  , .DOADO(
   {  r1do_31_, r1do_30_, r1do_29_, r1do_28_
  , r1do_27_, r1do_26_, r1do_25_, r1do_24_
  , r1do_23_, r1do_22_, r1do_21_, r1do_20_
  , r1do_19_, r1do_18_, r1do_17_, r1do_16_
  , r1do_15_, r1do_14_, r1do_13_, r1do_12_
  , r1do_11_, r1do_10_, r1do_9_, r1do_8_
  , r1do_7_, r1do_6_, r1do_5_, r1do_4_
  , r1do_3_, r1do_2_, r1do_1_, r1do_0_
   } )
  , .DOBDO(
   {  zsimv_ucon_29, zsimv_ucon_28, zsimv_ucon_26, zsimv_ucon_25
  , zsimv_ucon_24, zsimv_ucon_23, zsimv_ucon_22, zsimv_ucon_21
  , zsimv_ucon_20, zsimv_ucon_19, zsimv_ucon_18, zsimv_ucon_17
  , zsimv_ucon_15, zsimv_ucon_14, zsimv_ucon_13, zsimv_ucon_12
  , zsimv_ucon_11, zsimv_ucon_10, zsimv_ucon_9, zsimv_ucon_8
  , zsimv_ucon_7, zsimv_ucon_6, zsimv_ucon_36, zsimv_ucon_35
  , zsimv_ucon_34, zsimv_ucon_33, zsimv_ucon_32, zsimv_ucon_31
  , zsimv_ucon_30, zsimv_ucon_27, zsimv_ucon_16, RAMB36E1_DOBDO_0_
   } )
  );

defparam I_RAMB36E1_0.SRVAL_A = "000000000000000000000000000000000000";
defparam I_RAMB36E1_0.SRVAL_B = "000000000000000000000000000000000000";
defparam I_RAMB36E1_0.WRITE_MODE_A = "READ_FIRST";
defparam I_RAMB36E1_0.WRITE_MODE_B = "READ_FIRST";
defparam I_RAMB36E1_0.WRITE_WIDTH_B = 36;
defparam I_RAMB36E1_0.READ_WIDTH_A = 36;
RAMB36E1 I_RAMB36E1_0 (
    .CASCADEOUTA(zsimv_ucon_63)
  , .CASCADEOUTB(zsimv_ucon_64)
  , .DBITERR(zsimv_ucon_65)
  , .SBITERR(zsimv_ucon_118)
  , .CASCADEINA(zsimv_ucon_119)
  , .CASCADEINB(zsimv_ucon_120)
  , .CLKARDCLK(wire_sysFreq)
  , .CLKBWRCLK(w0clk)
  , .ENARDEN(alb_mss_mem_lat_0000_ZMEM_i_rdel_mem_add_vcc)
  , .ENBWREN(alb_mss_mem_lat_0000_ZMEM_i_rdel_mem_add_vcc)
  , .INJECTDBITERR(zsimv_ucon_121)
  , .INJECTSBITERR(zsimv_ucon_122)
  , .REGCEAREGCE(alb_mss_mem_lat_0000_ZMEM_i_rdel_mem_add_gnd)
  , .REGCEB(alb_mss_mem_lat_0000_ZMEM_i_rdel_mem_add_gnd)
  , .RSTRAMARSTRAM(alb_mss_mem_lat_0000_ZMEM_i_rdel_mem_add_gnd)
  , .RSTRAMB(alb_mss_mem_lat_0000_ZMEM_i_rdel_mem_add_gnd)
  , .RSTREGARSTREG(alb_mss_mem_lat_0000_ZMEM_i_rdel_mem_add_gnd)
  , .RSTREGB(alb_mss_mem_lat_0000_ZMEM_i_rdel_mem_add_gnd)
  , .DIPADIP(
   {  alb_mss_mem_lat_0000_ZMEM_i_rdel_mem_add_gnd, alb_mss_mem_lat_0000_ZMEM_i_rdel_mem_add_gnd, alb_mss_mem_lat_0000_ZMEM_i_rdel_mem_add_gnd, alb_mss_mem_lat_0000_ZMEM_i_rdel_mem_add_gnd
   } )
  , .DIPBDIP(
   {  w0di_71_, w0di_70_, w0di_69_, w0di_68_
   } )
  , .WEA(
   {  alb_mss_mem_lat_0000_ZMEM_i_rdel_mem_add_gnd, alb_mss_mem_lat_0000_ZMEM_i_rdel_mem_add_gnd, alb_mss_mem_lat_0000_ZMEM_i_rdel_mem_add_gnd, alb_mss_mem_lat_0000_ZMEM_i_rdel_mem_add_gnd
   } )
  , .WEBWE(
   {  w0we, w0we, w0we, w0we
  , w0we, w0we, w0we, w0we
   } )
  , .ADDRARDADDR(
   {  alb_mss_mem_lat_0000_ZMEM_i_rdel_mem_add_gnd, PROTECTED_SETUP_r1addr_9_, PROTECTED_SETUP_r1addr_8_, PROTECTED_SETUP_r1addr_7_
  , PROTECTED_SETUP_r1addr_6_, PROTECTED_SETUP_r1addr_5_, PROTECTED_SETUP_r1addr_4_, PROTECTED_SETUP_r1addr_3_
  , PROTECTED_SETUP_r1addr_2_, PROTECTED_SETUP_r1addr_1_, PROTECTED_SETUP_r1addr_0_, alb_mss_mem_lat_0000_ZMEM_i_rdel_mem_add_gnd
  , alb_mss_mem_lat_0000_ZMEM_i_rdel_mem_add_gnd, alb_mss_mem_lat_0000_ZMEM_i_rdel_mem_add_gnd, alb_mss_mem_lat_0000_ZMEM_i_rdel_mem_add_gnd, alb_mss_mem_lat_0000_ZMEM_i_rdel_mem_add_gnd
   } )
  , .ADDRBWRADDR(
   {  alb_mss_mem_lat_0000_ZMEM_i_rdel_mem_add_gnd, w0addr_9_, w0addr_8_, w0addr_7_
  , w0addr_6_, w0addr_5_, w0addr_4_, w0addr_3_
  , w0addr_2_, w0addr_1_, w0addr_0_, alb_mss_mem_lat_0000_ZMEM_i_rdel_mem_add_gnd
  , alb_mss_mem_lat_0000_ZMEM_i_rdel_mem_add_gnd, alb_mss_mem_lat_0000_ZMEM_i_rdel_mem_add_gnd, alb_mss_mem_lat_0000_ZMEM_i_rdel_mem_add_gnd, alb_mss_mem_lat_0000_ZMEM_i_rdel_mem_add_gnd
   } )
  , .DIADI(
   {  alb_mss_mem_lat_0000_ZMEM_i_rdel_mem_add_gnd, alb_mss_mem_lat_0000_ZMEM_i_rdel_mem_add_gnd, alb_mss_mem_lat_0000_ZMEM_i_rdel_mem_add_gnd, alb_mss_mem_lat_0000_ZMEM_i_rdel_mem_add_gnd
  , alb_mss_mem_lat_0000_ZMEM_i_rdel_mem_add_gnd, alb_mss_mem_lat_0000_ZMEM_i_rdel_mem_add_gnd, alb_mss_mem_lat_0000_ZMEM_i_rdel_mem_add_gnd, alb_mss_mem_lat_0000_ZMEM_i_rdel_mem_add_gnd
  , alb_mss_mem_lat_0000_ZMEM_i_rdel_mem_add_gnd, alb_mss_mem_lat_0000_ZMEM_i_rdel_mem_add_gnd, alb_mss_mem_lat_0000_ZMEM_i_rdel_mem_add_gnd, alb_mss_mem_lat_0000_ZMEM_i_rdel_mem_add_gnd
  , alb_mss_mem_lat_0000_ZMEM_i_rdel_mem_add_gnd, alb_mss_mem_lat_0000_ZMEM_i_rdel_mem_add_gnd, alb_mss_mem_lat_0000_ZMEM_i_rdel_mem_add_gnd, alb_mss_mem_lat_0000_ZMEM_i_rdel_mem_add_gnd
  , alb_mss_mem_lat_0000_ZMEM_i_rdel_mem_add_gnd, alb_mss_mem_lat_0000_ZMEM_i_rdel_mem_add_gnd, alb_mss_mem_lat_0000_ZMEM_i_rdel_mem_add_gnd, alb_mss_mem_lat_0000_ZMEM_i_rdel_mem_add_gnd
  , alb_mss_mem_lat_0000_ZMEM_i_rdel_mem_add_gnd, alb_mss_mem_lat_0000_ZMEM_i_rdel_mem_add_gnd, alb_mss_mem_lat_0000_ZMEM_i_rdel_mem_add_gnd, alb_mss_mem_lat_0000_ZMEM_i_rdel_mem_add_gnd
  , alb_mss_mem_lat_0000_ZMEM_i_rdel_mem_add_gnd, alb_mss_mem_lat_0000_ZMEM_i_rdel_mem_add_gnd, alb_mss_mem_lat_0000_ZMEM_i_rdel_mem_add_gnd, alb_mss_mem_lat_0000_ZMEM_i_rdel_mem_add_gnd
  , alb_mss_mem_lat_0000_ZMEM_i_rdel_mem_add_gnd, alb_mss_mem_lat_0000_ZMEM_i_rdel_mem_add_gnd, alb_mss_mem_lat_0000_ZMEM_i_rdel_mem_add_gnd, alb_mss_mem_lat_0000_ZMEM_i_rdel_mem_add_gnd
   } )
  , .DIBDI(
   {  w0di_67_, w0di_66_, w0di_65_, w0di_64_
  , w0di_63_, w0di_62_, w0di_61_, w0di_60_
  , w0di_59_, w0di_58_, w0di_57_, w0di_56_
  , w0di_55_, w0di_54_, w0di_53_, w0di_52_
  , w0di_51_, w0di_50_, w0di_49_, w0di_48_
  , w0di_47_, w0di_46_, w0di_45_, w0di_44_
  , w0di_43_, w0di_42_, w0di_41_, w0di_40_
  , w0di_39_, w0di_38_, w0di_37_, w0di_36_
   } )
  , .DOPADOP(
   {  r1do_71_, r1do_70_, r1do_69_, r1do_68_
   } )
  , .DOPBDOP(
   {  zsimv_ucon_100, zsimv_ucon_99, zsimv_ucon_98, zsimv_ucon_97
   } )
  , .ECCPARITY(
   {  zsimv_ucon_108, zsimv_ucon_107, zsimv_ucon_106, zsimv_ucon_105
  , zsimv_ucon_104, zsimv_ucon_103, zsimv_ucon_102, zsimv_ucon_101
   } )
  , .RDADDRECC(
   {  zsimv_ucon_117, zsimv_ucon_116, zsimv_ucon_115, zsimv_ucon_114
  , zsimv_ucon_113, zsimv_ucon_112, zsimv_ucon_111, zsimv_ucon_110
  , zsimv_ucon_109 } )
  , .DOADO(
   {  r1do_67_, r1do_66_, r1do_65_, r1do_64_
  , r1do_63_, r1do_62_, r1do_61_, r1do_60_
  , r1do_59_, r1do_58_, r1do_57_, r1do_56_
  , r1do_55_, r1do_54_, r1do_53_, r1do_52_
  , r1do_51_, r1do_50_, r1do_49_, r1do_48_
  , r1do_47_, r1do_46_, r1do_45_, r1do_44_
  , r1do_43_, r1do_42_, r1do_41_, r1do_40_
  , r1do_39_, r1do_38_, r1do_37_, r1do_36_
   } )
  , .DOBDO(
   {  zsimv_ucon_89, zsimv_ucon_88, zsimv_ucon_86, zsimv_ucon_85
  , zsimv_ucon_84, zsimv_ucon_83, zsimv_ucon_82, zsimv_ucon_81
  , zsimv_ucon_80, zsimv_ucon_79, zsimv_ucon_78, zsimv_ucon_77
  , zsimv_ucon_75, zsimv_ucon_74, zsimv_ucon_73, zsimv_ucon_72
  , zsimv_ucon_71, zsimv_ucon_70, zsimv_ucon_69, zsimv_ucon_68
  , zsimv_ucon_67, zsimv_ucon_66, zsimv_ucon_96, zsimv_ucon_95
  , zsimv_ucon_94, zsimv_ucon_93, zsimv_ucon_92, zsimv_ucon_91
  , zsimv_ucon_90, zsimv_ucon_87, zsimv_ucon_76, RAMB36E1_0_DOBDO_0_
   } )
  );

defparam I_RAMB36E1_1.SRVAL_A = "000000000000000000000000000000000000";
defparam I_RAMB36E1_1.SRVAL_B = "000000000000000000000000000000000000";
defparam I_RAMB36E1_1.WRITE_MODE_A = "READ_FIRST";
defparam I_RAMB36E1_1.WRITE_MODE_B = "READ_FIRST";
defparam I_RAMB36E1_1.WRITE_WIDTH_B = 36;
defparam I_RAMB36E1_1.READ_WIDTH_A = 36;
RAMB36E1 I_RAMB36E1_1 (
    .CASCADEOUTA(zsimv_ucon_123)
  , .CASCADEOUTB(zsimv_ucon_124)
  , .DBITERR(zsimv_ucon_125)
  , .SBITERR(zsimv_ucon_178)
  , .CASCADEINA(zsimv_ucon_179)
  , .CASCADEINB(zsimv_ucon_180)
  , .CLKARDCLK(wire_sysFreq)
  , .CLKBWRCLK(w0clk)
  , .ENARDEN(alb_mss_mem_lat_0000_ZMEM_i_rdel_mem_add_vcc)
  , .ENBWREN(alb_mss_mem_lat_0000_ZMEM_i_rdel_mem_add_vcc)
  , .INJECTDBITERR(zsimv_ucon_181)
  , .INJECTSBITERR(zsimv_ucon_182)
  , .REGCEAREGCE(alb_mss_mem_lat_0000_ZMEM_i_rdel_mem_add_gnd)
  , .REGCEB(alb_mss_mem_lat_0000_ZMEM_i_rdel_mem_add_gnd)
  , .RSTRAMARSTRAM(alb_mss_mem_lat_0000_ZMEM_i_rdel_mem_add_gnd)
  , .RSTRAMB(alb_mss_mem_lat_0000_ZMEM_i_rdel_mem_add_gnd)
  , .RSTREGARSTREG(alb_mss_mem_lat_0000_ZMEM_i_rdel_mem_add_gnd)
  , .RSTREGB(alb_mss_mem_lat_0000_ZMEM_i_rdel_mem_add_gnd)
  , .DIPADIP(
   {  alb_mss_mem_lat_0000_ZMEM_i_rdel_mem_add_gnd, alb_mss_mem_lat_0000_ZMEM_i_rdel_mem_add_gnd, alb_mss_mem_lat_0000_ZMEM_i_rdel_mem_add_gnd, alb_mss_mem_lat_0000_ZMEM_i_rdel_mem_add_gnd
   } )
  , .DIPBDIP(
   {  w0di_107_, w0di_106_, w0di_105_, w0di_104_
   } )
  , .WEA(
   {  alb_mss_mem_lat_0000_ZMEM_i_rdel_mem_add_gnd, alb_mss_mem_lat_0000_ZMEM_i_rdel_mem_add_gnd, alb_mss_mem_lat_0000_ZMEM_i_rdel_mem_add_gnd, alb_mss_mem_lat_0000_ZMEM_i_rdel_mem_add_gnd
   } )
  , .WEBWE(
   {  w0we, w0we, w0we, w0we
  , w0we, w0we, w0we, w0we
   } )
  , .ADDRARDADDR(
   {  alb_mss_mem_lat_0000_ZMEM_i_rdel_mem_add_gnd, PROTECTED_SETUP_r1addr_9_, PROTECTED_SETUP_r1addr_8_, PROTECTED_SETUP_r1addr_7_
  , PROTECTED_SETUP_r1addr_6_, PROTECTED_SETUP_r1addr_5_, PROTECTED_SETUP_r1addr_4_, PROTECTED_SETUP_r1addr_3_
  , PROTECTED_SETUP_r1addr_2_, PROTECTED_SETUP_r1addr_1_, PROTECTED_SETUP_r1addr_0_, alb_mss_mem_lat_0000_ZMEM_i_rdel_mem_add_gnd
  , alb_mss_mem_lat_0000_ZMEM_i_rdel_mem_add_gnd, alb_mss_mem_lat_0000_ZMEM_i_rdel_mem_add_gnd, alb_mss_mem_lat_0000_ZMEM_i_rdel_mem_add_gnd, alb_mss_mem_lat_0000_ZMEM_i_rdel_mem_add_gnd
   } )
  , .ADDRBWRADDR(
   {  alb_mss_mem_lat_0000_ZMEM_i_rdel_mem_add_gnd, w0addr_9_, w0addr_8_, w0addr_7_
  , w0addr_6_, w0addr_5_, w0addr_4_, w0addr_3_
  , w0addr_2_, w0addr_1_, w0addr_0_, alb_mss_mem_lat_0000_ZMEM_i_rdel_mem_add_gnd
  , alb_mss_mem_lat_0000_ZMEM_i_rdel_mem_add_gnd, alb_mss_mem_lat_0000_ZMEM_i_rdel_mem_add_gnd, alb_mss_mem_lat_0000_ZMEM_i_rdel_mem_add_gnd, alb_mss_mem_lat_0000_ZMEM_i_rdel_mem_add_gnd
   } )
  , .DIADI(
   {  alb_mss_mem_lat_0000_ZMEM_i_rdel_mem_add_gnd, alb_mss_mem_lat_0000_ZMEM_i_rdel_mem_add_gnd, alb_mss_mem_lat_0000_ZMEM_i_rdel_mem_add_gnd, alb_mss_mem_lat_0000_ZMEM_i_rdel_mem_add_gnd
  , alb_mss_mem_lat_0000_ZMEM_i_rdel_mem_add_gnd, alb_mss_mem_lat_0000_ZMEM_i_rdel_mem_add_gnd, alb_mss_mem_lat_0000_ZMEM_i_rdel_mem_add_gnd, alb_mss_mem_lat_0000_ZMEM_i_rdel_mem_add_gnd
  , alb_mss_mem_lat_0000_ZMEM_i_rdel_mem_add_gnd, alb_mss_mem_lat_0000_ZMEM_i_rdel_mem_add_gnd, alb_mss_mem_lat_0000_ZMEM_i_rdel_mem_add_gnd, alb_mss_mem_lat_0000_ZMEM_i_rdel_mem_add_gnd
  , alb_mss_mem_lat_0000_ZMEM_i_rdel_mem_add_gnd, alb_mss_mem_lat_0000_ZMEM_i_rdel_mem_add_gnd, alb_mss_mem_lat_0000_ZMEM_i_rdel_mem_add_gnd, alb_mss_mem_lat_0000_ZMEM_i_rdel_mem_add_gnd
  , alb_mss_mem_lat_0000_ZMEM_i_rdel_mem_add_gnd, alb_mss_mem_lat_0000_ZMEM_i_rdel_mem_add_gnd, alb_mss_mem_lat_0000_ZMEM_i_rdel_mem_add_gnd, alb_mss_mem_lat_0000_ZMEM_i_rdel_mem_add_gnd
  , alb_mss_mem_lat_0000_ZMEM_i_rdel_mem_add_gnd, alb_mss_mem_lat_0000_ZMEM_i_rdel_mem_add_gnd, alb_mss_mem_lat_0000_ZMEM_i_rdel_mem_add_gnd, alb_mss_mem_lat_0000_ZMEM_i_rdel_mem_add_gnd
  , alb_mss_mem_lat_0000_ZMEM_i_rdel_mem_add_gnd, alb_mss_mem_lat_0000_ZMEM_i_rdel_mem_add_gnd, alb_mss_mem_lat_0000_ZMEM_i_rdel_mem_add_gnd, alb_mss_mem_lat_0000_ZMEM_i_rdel_mem_add_gnd
  , alb_mss_mem_lat_0000_ZMEM_i_rdel_mem_add_gnd, alb_mss_mem_lat_0000_ZMEM_i_rdel_mem_add_gnd, alb_mss_mem_lat_0000_ZMEM_i_rdel_mem_add_gnd, alb_mss_mem_lat_0000_ZMEM_i_rdel_mem_add_gnd
   } )
  , .DIBDI(
   {  w0di_103_, w0di_102_, w0di_101_, w0di_100_
  , w0di_99_, w0di_98_, w0di_97_, w0di_96_
  , w0di_95_, w0di_94_, w0di_93_, w0di_92_
  , w0di_91_, w0di_90_, w0di_89_, w0di_88_
  , w0di_87_, w0di_86_, w0di_85_, w0di_84_
  , w0di_83_, w0di_82_, w0di_81_, w0di_80_
  , w0di_79_, w0di_78_, w0di_77_, w0di_76_
  , w0di_75_, w0di_74_, w0di_73_, w0di_72_
   } )
  , .DOPADOP(
   {  r1do_107_, r1do_106_, r1do_105_, r1do_104_
   } )
  , .DOPBDOP(
   {  zsimv_ucon_160, zsimv_ucon_159, zsimv_ucon_158, zsimv_ucon_157
   } )
  , .ECCPARITY(
   {  zsimv_ucon_168, zsimv_ucon_167, zsimv_ucon_166, zsimv_ucon_165
  , zsimv_ucon_164, zsimv_ucon_163, zsimv_ucon_162, zsimv_ucon_161
   } )
  , .RDADDRECC(
   {  zsimv_ucon_177, zsimv_ucon_176, zsimv_ucon_175, zsimv_ucon_174
  , zsimv_ucon_173, zsimv_ucon_172, zsimv_ucon_171, zsimv_ucon_170
  , zsimv_ucon_169 } )
  , .DOADO(
   {  r1do_103_, r1do_102_, r1do_101_, r1do_100_
  , r1do_99_, r1do_98_, r1do_97_, r1do_96_
  , r1do_95_, r1do_94_, r1do_93_, r1do_92_
  , r1do_91_, r1do_90_, r1do_89_, r1do_88_
  , r1do_87_, r1do_86_, r1do_85_, r1do_84_
  , r1do_83_, r1do_82_, r1do_81_, r1do_80_
  , r1do_79_, r1do_78_, r1do_77_, r1do_76_
  , r1do_75_, r1do_74_, r1do_73_, r1do_72_
   } )
  , .DOBDO(
   {  zsimv_ucon_149, zsimv_ucon_148, zsimv_ucon_146, zsimv_ucon_145
  , zsimv_ucon_144, zsimv_ucon_143, zsimv_ucon_142, zsimv_ucon_141
  , zsimv_ucon_140, zsimv_ucon_139, zsimv_ucon_138, zsimv_ucon_137
  , zsimv_ucon_135, zsimv_ucon_134, zsimv_ucon_133, zsimv_ucon_132
  , zsimv_ucon_131, zsimv_ucon_130, zsimv_ucon_129, zsimv_ucon_128
  , zsimv_ucon_127, zsimv_ucon_126, zsimv_ucon_156, zsimv_ucon_155
  , zsimv_ucon_154, zsimv_ucon_153, zsimv_ucon_152, zsimv_ucon_151
  , zsimv_ucon_150, zsimv_ucon_147, zsimv_ucon_136, RAMB36E1_1_DOBDO_0_
   } )
  );

defparam I_RAMB36E1_2.SRVAL_A = "000000000000000000000000000000000000";
defparam I_RAMB36E1_2.SRVAL_B = "000000000000000000000000000000000000";
defparam I_RAMB36E1_2.WRITE_MODE_A = "READ_FIRST";
defparam I_RAMB36E1_2.WRITE_MODE_B = "READ_FIRST";
defparam I_RAMB36E1_2.WRITE_WIDTH_B = 36;
defparam I_RAMB36E1_2.READ_WIDTH_A = 36;
RAMB36E1 I_RAMB36E1_2 (
    .CASCADEOUTA(zsimv_ucon_183)
  , .CASCADEOUTB(zsimv_ucon_184)
  , .DBITERR(zsimv_ucon_185)
  , .SBITERR(zsimv_ucon_251)
  , .CASCADEINA(zsimv_ucon_252)
  , .CASCADEINB(zsimv_ucon_253)
  , .CLKARDCLK(wire_sysFreq)
  , .CLKBWRCLK(w0clk)
  , .ENARDEN(alb_mss_mem_lat_0000_ZMEM_i_rdel_mem_add_vcc)
  , .ENBWREN(alb_mss_mem_lat_0000_ZMEM_i_rdel_mem_add_vcc)
  , .INJECTDBITERR(zsimv_ucon_254)
  , .INJECTSBITERR(zsimv_ucon_255)
  , .REGCEAREGCE(alb_mss_mem_lat_0000_ZMEM_i_rdel_mem_add_gnd)
  , .REGCEB(alb_mss_mem_lat_0000_ZMEM_i_rdel_mem_add_gnd)
  , .RSTRAMARSTRAM(alb_mss_mem_lat_0000_ZMEM_i_rdel_mem_add_gnd)
  , .RSTRAMB(alb_mss_mem_lat_0000_ZMEM_i_rdel_mem_add_gnd)
  , .RSTREGARSTREG(alb_mss_mem_lat_0000_ZMEM_i_rdel_mem_add_gnd)
  , .RSTREGB(alb_mss_mem_lat_0000_ZMEM_i_rdel_mem_add_gnd)
  , .DIPADIP(
   {  alb_mss_mem_lat_0000_ZMEM_i_rdel_mem_add_gnd, alb_mss_mem_lat_0000_ZMEM_i_rdel_mem_add_gnd, alb_mss_mem_lat_0000_ZMEM_i_rdel_mem_add_gnd, alb_mss_mem_lat_0000_ZMEM_i_rdel_mem_add_gnd
   } )
  , .DIPBDIP(
   {  alb_mss_mem_lat_0000_ZMEM_i_rdel_mem_add_gnd, alb_mss_mem_lat_0000_ZMEM_i_rdel_mem_add_gnd, alb_mss_mem_lat_0000_ZMEM_i_rdel_mem_add_gnd, alb_mss_mem_lat_0000_ZMEM_i_rdel_mem_add_gnd
   } )
  , .WEA(
   {  alb_mss_mem_lat_0000_ZMEM_i_rdel_mem_add_gnd, alb_mss_mem_lat_0000_ZMEM_i_rdel_mem_add_gnd, alb_mss_mem_lat_0000_ZMEM_i_rdel_mem_add_gnd, alb_mss_mem_lat_0000_ZMEM_i_rdel_mem_add_gnd
   } )
  , .WEBWE(
   {  w0we, w0we, w0we, w0we
  , w0we, w0we, w0we, w0we
   } )
  , .ADDRARDADDR(
   {  alb_mss_mem_lat_0000_ZMEM_i_rdel_mem_add_gnd, PROTECTED_SETUP_r1addr_9_, PROTECTED_SETUP_r1addr_8_, PROTECTED_SETUP_r1addr_7_
  , PROTECTED_SETUP_r1addr_6_, PROTECTED_SETUP_r1addr_5_, PROTECTED_SETUP_r1addr_4_, PROTECTED_SETUP_r1addr_3_
  , PROTECTED_SETUP_r1addr_2_, PROTECTED_SETUP_r1addr_1_, PROTECTED_SETUP_r1addr_0_, alb_mss_mem_lat_0000_ZMEM_i_rdel_mem_add_gnd
  , alb_mss_mem_lat_0000_ZMEM_i_rdel_mem_add_gnd, alb_mss_mem_lat_0000_ZMEM_i_rdel_mem_add_gnd, alb_mss_mem_lat_0000_ZMEM_i_rdel_mem_add_gnd, alb_mss_mem_lat_0000_ZMEM_i_rdel_mem_add_gnd
   } )
  , .ADDRBWRADDR(
   {  alb_mss_mem_lat_0000_ZMEM_i_rdel_mem_add_gnd, w0addr_9_, w0addr_8_, w0addr_7_
  , w0addr_6_, w0addr_5_, w0addr_4_, w0addr_3_
  , w0addr_2_, w0addr_1_, w0addr_0_, alb_mss_mem_lat_0000_ZMEM_i_rdel_mem_add_gnd
  , alb_mss_mem_lat_0000_ZMEM_i_rdel_mem_add_gnd, alb_mss_mem_lat_0000_ZMEM_i_rdel_mem_add_gnd, alb_mss_mem_lat_0000_ZMEM_i_rdel_mem_add_gnd, alb_mss_mem_lat_0000_ZMEM_i_rdel_mem_add_gnd
   } )
  , .DIADI(
   {  alb_mss_mem_lat_0000_ZMEM_i_rdel_mem_add_gnd, alb_mss_mem_lat_0000_ZMEM_i_rdel_mem_add_gnd, alb_mss_mem_lat_0000_ZMEM_i_rdel_mem_add_gnd, alb_mss_mem_lat_0000_ZMEM_i_rdel_mem_add_gnd
  , alb_mss_mem_lat_0000_ZMEM_i_rdel_mem_add_gnd, alb_mss_mem_lat_0000_ZMEM_i_rdel_mem_add_gnd, alb_mss_mem_lat_0000_ZMEM_i_rdel_mem_add_gnd, alb_mss_mem_lat_0000_ZMEM_i_rdel_mem_add_gnd
  , alb_mss_mem_lat_0000_ZMEM_i_rdel_mem_add_gnd, alb_mss_mem_lat_0000_ZMEM_i_rdel_mem_add_gnd, alb_mss_mem_lat_0000_ZMEM_i_rdel_mem_add_gnd, alb_mss_mem_lat_0000_ZMEM_i_rdel_mem_add_gnd
  , alb_mss_mem_lat_0000_ZMEM_i_rdel_mem_add_gnd, alb_mss_mem_lat_0000_ZMEM_i_rdel_mem_add_gnd, alb_mss_mem_lat_0000_ZMEM_i_rdel_mem_add_gnd, alb_mss_mem_lat_0000_ZMEM_i_rdel_mem_add_gnd
  , alb_mss_mem_lat_0000_ZMEM_i_rdel_mem_add_gnd, alb_mss_mem_lat_0000_ZMEM_i_rdel_mem_add_gnd, alb_mss_mem_lat_0000_ZMEM_i_rdel_mem_add_gnd, alb_mss_mem_lat_0000_ZMEM_i_rdel_mem_add_gnd
  , alb_mss_mem_lat_0000_ZMEM_i_rdel_mem_add_gnd, alb_mss_mem_lat_0000_ZMEM_i_rdel_mem_add_gnd, alb_mss_mem_lat_0000_ZMEM_i_rdel_mem_add_gnd, alb_mss_mem_lat_0000_ZMEM_i_rdel_mem_add_gnd
  , alb_mss_mem_lat_0000_ZMEM_i_rdel_mem_add_gnd, alb_mss_mem_lat_0000_ZMEM_i_rdel_mem_add_gnd, alb_mss_mem_lat_0000_ZMEM_i_rdel_mem_add_gnd, alb_mss_mem_lat_0000_ZMEM_i_rdel_mem_add_gnd
  , alb_mss_mem_lat_0000_ZMEM_i_rdel_mem_add_gnd, alb_mss_mem_lat_0000_ZMEM_i_rdel_mem_add_gnd, alb_mss_mem_lat_0000_ZMEM_i_rdel_mem_add_gnd, alb_mss_mem_lat_0000_ZMEM_i_rdel_mem_add_gnd
   } )
  , .DIBDI(
   {  alb_mss_mem_lat_0000_ZMEM_i_rdel_mem_add_gnd, alb_mss_mem_lat_0000_ZMEM_i_rdel_mem_add_gnd, alb_mss_mem_lat_0000_ZMEM_i_rdel_mem_add_gnd, alb_mss_mem_lat_0000_ZMEM_i_rdel_mem_add_gnd
  , alb_mss_mem_lat_0000_ZMEM_i_rdel_mem_add_gnd, alb_mss_mem_lat_0000_ZMEM_i_rdel_mem_add_gnd, alb_mss_mem_lat_0000_ZMEM_i_rdel_mem_add_gnd, alb_mss_mem_lat_0000_ZMEM_i_rdel_mem_add_gnd
  , alb_mss_mem_lat_0000_ZMEM_i_rdel_mem_add_gnd, w0di_130_, w0di_129_, w0di_128_
  , w0di_127_, w0di_126_, w0di_125_, w0di_124_
  , w0di_123_, w0di_122_, w0di_121_, w0di_120_
  , w0di_119_, w0di_118_, w0di_117_, w0di_116_
  , w0di_115_, w0di_114_, w0di_113_, w0di_112_
  , w0di_111_, w0di_110_, w0di_109_, w0di_108_
   } )
  , .DOPADOP(
   {  zsimv_ucon_229, zsimv_ucon_228, zsimv_ucon_227, zsimv_ucon_226
   } )
  , .DOPBDOP(
   {  zsimv_ucon_233, zsimv_ucon_232, zsimv_ucon_231, zsimv_ucon_230
   } )
  , .ECCPARITY(
   {  zsimv_ucon_241, zsimv_ucon_240, zsimv_ucon_239, zsimv_ucon_238
  , zsimv_ucon_237, zsimv_ucon_236, zsimv_ucon_235, zsimv_ucon_234
   } )
  , .RDADDRECC(
   {  zsimv_ucon_250, zsimv_ucon_249, zsimv_ucon_248, zsimv_ucon_247
  , zsimv_ucon_246, zsimv_ucon_245, zsimv_ucon_244, zsimv_ucon_243
  , zsimv_ucon_242 } )
  , .DOADO(
   {  zsimv_ucon_194, zsimv_ucon_193, zsimv_ucon_192, zsimv_ucon_191
  , zsimv_ucon_190, zsimv_ucon_189, zsimv_ucon_188, zsimv_ucon_187
  , zsimv_ucon_186, r1do_130_, r1do_129_, r1do_128_
  , r1do_127_, r1do_126_, r1do_125_, r1do_124_
  , r1do_123_, r1do_122_, r1do_121_, r1do_120_
  , r1do_119_, r1do_118_, r1do_117_, r1do_116_
  , r1do_115_, r1do_114_, r1do_113_, r1do_112_
  , r1do_111_, r1do_110_, r1do_109_, r1do_108_
   } )
  , .DOBDO(
   {  zsimv_ucon_218, zsimv_ucon_217, zsimv_ucon_215, zsimv_ucon_214
  , zsimv_ucon_213, zsimv_ucon_212, zsimv_ucon_211, zsimv_ucon_210
  , zsimv_ucon_209, zsimv_ucon_208, zsimv_ucon_207, zsimv_ucon_206
  , zsimv_ucon_204, zsimv_ucon_203, zsimv_ucon_202, zsimv_ucon_201
  , zsimv_ucon_200, zsimv_ucon_199, zsimv_ucon_198, zsimv_ucon_197
  , zsimv_ucon_196, zsimv_ucon_195, zsimv_ucon_225, zsimv_ucon_224
  , zsimv_ucon_223, zsimv_ucon_222, zsimv_ucon_221, zsimv_ucon_220
  , zsimv_ucon_219, zsimv_ucon_216, zsimv_ucon_205, RAMB36E1_2_DOBDO_0_
   } )
  );

zview I_zview_w0we (
    .I(w0we)
  );

zview \I_zview_w0addr[9]  (
    .I(w0addr_9_)
  );

zview \I_zview_w0addr[8]  (
    .I(w0addr_8_)
  );

zview \I_zview_w0addr[7]  (
    .I(w0addr_7_)
  );

zview \I_zview_w0addr[6]  (
    .I(w0addr_6_)
  );

zview \I_zview_w0addr[5]  (
    .I(w0addr_5_)
  );

zview \I_zview_w0addr[4]  (
    .I(w0addr_4_)
  );

zview \I_zview_w0addr[3]  (
    .I(w0addr_3_)
  );

zview \I_zview_w0addr[2]  (
    .I(w0addr_2_)
  );

zview \I_zview_w0addr[1]  (
    .I(w0addr_1_)
  );

zview \I_zview_w0addr[0]  (
    .I(w0addr_0_)
  );

zview \I_zview_w0di[130]  (
    .I(w0di_130_)
  );

zview \I_zview_w0di[129]  (
    .I(w0di_129_)
  );

zview \I_zview_w0di[128]  (
    .I(w0di_128_)
  );

zview \I_zview_w0di[127]  (
    .I(w0di_127_)
  );

zview \I_zview_w0di[126]  (
    .I(w0di_126_)
  );

zview \I_zview_w0di[125]  (
    .I(w0di_125_)
  );

zview \I_zview_w0di[124]  (
    .I(w0di_124_)
  );

zview \I_zview_w0di[123]  (
    .I(w0di_123_)
  );

zview \I_zview_w0di[122]  (
    .I(w0di_122_)
  );

zview \I_zview_w0di[121]  (
    .I(w0di_121_)
  );

zview \I_zview_w0di[120]  (
    .I(w0di_120_)
  );

zview \I_zview_w0di[119]  (
    .I(w0di_119_)
  );

zview \I_zview_w0di[118]  (
    .I(w0di_118_)
  );

zview \I_zview_w0di[117]  (
    .I(w0di_117_)
  );

zview \I_zview_w0di[116]  (
    .I(w0di_116_)
  );

zview \I_zview_w0di[115]  (
    .I(w0di_115_)
  );

zview \I_zview_w0di[114]  (
    .I(w0di_114_)
  );

zview \I_zview_w0di[113]  (
    .I(w0di_113_)
  );

zview \I_zview_w0di[112]  (
    .I(w0di_112_)
  );

zview \I_zview_w0di[111]  (
    .I(w0di_111_)
  );

zview \I_zview_w0di[110]  (
    .I(w0di_110_)
  );

zview \I_zview_w0di[109]  (
    .I(w0di_109_)
  );

zview \I_zview_w0di[108]  (
    .I(w0di_108_)
  );

zview \I_zview_w0di[107]  (
    .I(w0di_107_)
  );

zview \I_zview_w0di[106]  (
    .I(w0di_106_)
  );

zview \I_zview_w0di[105]  (
    .I(w0di_105_)
  );

zview \I_zview_w0di[104]  (
    .I(w0di_104_)
  );

zview \I_zview_w0di[103]  (
    .I(w0di_103_)
  );

zview \I_zview_w0di[102]  (
    .I(w0di_102_)
  );

zview \I_zview_w0di[101]  (
    .I(w0di_101_)
  );

zview \I_zview_w0di[100]  (
    .I(w0di_100_)
  );

zview \I_zview_w0di[99]  (
    .I(w0di_99_)
  );

zview \I_zview_w0di[98]  (
    .I(w0di_98_)
  );

zview \I_zview_w0di[97]  (
    .I(w0di_97_)
  );

zview \I_zview_w0di[96]  (
    .I(w0di_96_)
  );

zview \I_zview_w0di[95]  (
    .I(w0di_95_)
  );

zview \I_zview_w0di[94]  (
    .I(w0di_94_)
  );

zview \I_zview_w0di[93]  (
    .I(w0di_93_)
  );

zview \I_zview_w0di[92]  (
    .I(w0di_92_)
  );

zview \I_zview_w0di[91]  (
    .I(w0di_91_)
  );

zview \I_zview_w0di[90]  (
    .I(w0di_90_)
  );

zview \I_zview_w0di[89]  (
    .I(w0di_89_)
  );

zview \I_zview_w0di[88]  (
    .I(w0di_88_)
  );

zview \I_zview_w0di[87]  (
    .I(w0di_87_)
  );

zview \I_zview_w0di[86]  (
    .I(w0di_86_)
  );

zview \I_zview_w0di[85]  (
    .I(w0di_85_)
  );

zview \I_zview_w0di[84]  (
    .I(w0di_84_)
  );

zview \I_zview_w0di[83]  (
    .I(w0di_83_)
  );

zview \I_zview_w0di[82]  (
    .I(w0di_82_)
  );

zview \I_zview_w0di[81]  (
    .I(w0di_81_)
  );

zview \I_zview_w0di[80]  (
    .I(w0di_80_)
  );

zview \I_zview_w0di[79]  (
    .I(w0di_79_)
  );

zview \I_zview_w0di[78]  (
    .I(w0di_78_)
  );

zview \I_zview_w0di[77]  (
    .I(w0di_77_)
  );

zview \I_zview_w0di[76]  (
    .I(w0di_76_)
  );

zview \I_zview_w0di[75]  (
    .I(w0di_75_)
  );

zview \I_zview_w0di[74]  (
    .I(w0di_74_)
  );

zview \I_zview_w0di[73]  (
    .I(w0di_73_)
  );

zview \I_zview_w0di[72]  (
    .I(w0di_72_)
  );

zview \I_zview_w0di[71]  (
    .I(w0di_71_)
  );

zview \I_zview_w0di[70]  (
    .I(w0di_70_)
  );

zview \I_zview_w0di[69]  (
    .I(w0di_69_)
  );

zview \I_zview_w0di[68]  (
    .I(w0di_68_)
  );

zview \I_zview_w0di[67]  (
    .I(w0di_67_)
  );

zview \I_zview_w0di[66]  (
    .I(w0di_66_)
  );

zview \I_zview_w0di[65]  (
    .I(w0di_65_)
  );

zview \I_zview_w0di[64]  (
    .I(w0di_64_)
  );

zview \I_zview_w0di[63]  (
    .I(w0di_63_)
  );

zview \I_zview_w0di[62]  (
    .I(w0di_62_)
  );

zview \I_zview_w0di[61]  (
    .I(w0di_61_)
  );

zview \I_zview_w0di[60]  (
    .I(w0di_60_)
  );

zview \I_zview_w0di[59]  (
    .I(w0di_59_)
  );

zview \I_zview_w0di[58]  (
    .I(w0di_58_)
  );

zview \I_zview_w0di[57]  (
    .I(w0di_57_)
  );

zview \I_zview_w0di[56]  (
    .I(w0di_56_)
  );

zview \I_zview_w0di[55]  (
    .I(w0di_55_)
  );

zview \I_zview_w0di[54]  (
    .I(w0di_54_)
  );

zview \I_zview_w0di[53]  (
    .I(w0di_53_)
  );

zview \I_zview_w0di[52]  (
    .I(w0di_52_)
  );

zview \I_zview_w0di[51]  (
    .I(w0di_51_)
  );

zview \I_zview_w0di[50]  (
    .I(w0di_50_)
  );

zview \I_zview_w0di[49]  (
    .I(w0di_49_)
  );

zview \I_zview_w0di[48]  (
    .I(w0di_48_)
  );

zview \I_zview_w0di[47]  (
    .I(w0di_47_)
  );

zview \I_zview_w0di[46]  (
    .I(w0di_46_)
  );

zview \I_zview_w0di[45]  (
    .I(w0di_45_)
  );

zview \I_zview_w0di[44]  (
    .I(w0di_44_)
  );

zview \I_zview_w0di[43]  (
    .I(w0di_43_)
  );

zview \I_zview_w0di[42]  (
    .I(w0di_42_)
  );

zview \I_zview_w0di[41]  (
    .I(w0di_41_)
  );

zview \I_zview_w0di[40]  (
    .I(w0di_40_)
  );

zview \I_zview_w0di[39]  (
    .I(w0di_39_)
  );

zview \I_zview_w0di[38]  (
    .I(w0di_38_)
  );

zview \I_zview_w0di[37]  (
    .I(w0di_37_)
  );

zview \I_zview_w0di[36]  (
    .I(w0di_36_)
  );

zview \I_zview_w0di[35]  (
    .I(w0di_35_)
  );

zview \I_zview_w0di[34]  (
    .I(w0di_34_)
  );

zview \I_zview_w0di[33]  (
    .I(w0di_33_)
  );

zview \I_zview_w0di[32]  (
    .I(w0di_32_)
  );

zview \I_zview_w0di[31]  (
    .I(w0di_31_)
  );

zview \I_zview_w0di[30]  (
    .I(w0di_30_)
  );

zview \I_zview_w0di[29]  (
    .I(w0di_29_)
  );

zview \I_zview_w0di[28]  (
    .I(w0di_28_)
  );

zview \I_zview_w0di[27]  (
    .I(w0di_27_)
  );

zview \I_zview_w0di[26]  (
    .I(w0di_26_)
  );

zview \I_zview_w0di[25]  (
    .I(w0di_25_)
  );

zview \I_zview_w0di[24]  (
    .I(w0di_24_)
  );

zview \I_zview_w0di[23]  (
    .I(w0di_23_)
  );

zview \I_zview_w0di[22]  (
    .I(w0di_22_)
  );

zview \I_zview_w0di[21]  (
    .I(w0di_21_)
  );

zview \I_zview_w0di[20]  (
    .I(w0di_20_)
  );

zview \I_zview_w0di[19]  (
    .I(w0di_19_)
  );

zview \I_zview_w0di[18]  (
    .I(w0di_18_)
  );

zview \I_zview_w0di[17]  (
    .I(w0di_17_)
  );

zview \I_zview_w0di[16]  (
    .I(w0di_16_)
  );

zview \I_zview_w0di[15]  (
    .I(w0di_15_)
  );

zview \I_zview_w0di[14]  (
    .I(w0di_14_)
  );

zview \I_zview_w0di[13]  (
    .I(w0di_13_)
  );

zview \I_zview_w0di[12]  (
    .I(w0di_12_)
  );

zview \I_zview_w0di[11]  (
    .I(w0di_11_)
  );

zview \I_zview_w0di[10]  (
    .I(w0di_10_)
  );

zview \I_zview_w0di[9]  (
    .I(w0di_9_)
  );

zview \I_zview_w0di[8]  (
    .I(w0di_8_)
  );

zview \I_zview_w0di[7]  (
    .I(w0di_7_)
  );

zview \I_zview_w0di[6]  (
    .I(w0di_6_)
  );

zview \I_zview_w0di[5]  (
    .I(w0di_5_)
  );

zview \I_zview_w0di[4]  (
    .I(w0di_4_)
  );

zview \I_zview_w0di[3]  (
    .I(w0di_3_)
  );

zview \I_zview_w0di[2]  (
    .I(w0di_2_)
  );

zview \I_zview_w0di[1]  (
    .I(w0di_1_)
  );

zview \I_zview_w0di[0]  (
    .I(w0di_0_)
  );

zview \I_zview_r1addr[9]  (
    .I(r1addr_9_)
  );

zview \I_zview_r1addr[8]  (
    .I(r1addr_8_)
  );

zview \I_zview_r1addr[7]  (
    .I(r1addr_7_)
  );

zview \I_zview_r1addr[6]  (
    .I(r1addr_6_)
  );

zview \I_zview_r1addr[5]  (
    .I(r1addr_5_)
  );

zview \I_zview_r1addr[4]  (
    .I(r1addr_4_)
  );

zview \I_zview_r1addr[3]  (
    .I(r1addr_3_)
  );

zview \I_zview_r1addr[2]  (
    .I(r1addr_2_)
  );

zview \I_zview_r1addr[1]  (
    .I(r1addr_1_)
  );

zview \I_zview_r1addr[0]  (
    .I(r1addr_0_)
  );

zview \I_zview_r1do[130]  (
    .I(r1do_130_)
  );

zview \I_zview_r1do[129]  (
    .I(r1do_129_)
  );

zview \I_zview_r1do[128]  (
    .I(r1do_128_)
  );

zview \I_zview_r1do[127]  (
    .I(r1do_127_)
  );

zview \I_zview_r1do[126]  (
    .I(r1do_126_)
  );

zview \I_zview_r1do[125]  (
    .I(r1do_125_)
  );

zview \I_zview_r1do[124]  (
    .I(r1do_124_)
  );

zview \I_zview_r1do[123]  (
    .I(r1do_123_)
  );

zview \I_zview_r1do[122]  (
    .I(r1do_122_)
  );

zview \I_zview_r1do[121]  (
    .I(r1do_121_)
  );

zview \I_zview_r1do[120]  (
    .I(r1do_120_)
  );

zview \I_zview_r1do[119]  (
    .I(r1do_119_)
  );

zview \I_zview_r1do[118]  (
    .I(r1do_118_)
  );

zview \I_zview_r1do[117]  (
    .I(r1do_117_)
  );

zview \I_zview_r1do[116]  (
    .I(r1do_116_)
  );

zview \I_zview_r1do[115]  (
    .I(r1do_115_)
  );

zview \I_zview_r1do[114]  (
    .I(r1do_114_)
  );

zview \I_zview_r1do[113]  (
    .I(r1do_113_)
  );

zview \I_zview_r1do[112]  (
    .I(r1do_112_)
  );

zview \I_zview_r1do[111]  (
    .I(r1do_111_)
  );

zview \I_zview_r1do[110]  (
    .I(r1do_110_)
  );

zview \I_zview_r1do[109]  (
    .I(r1do_109_)
  );

zview \I_zview_r1do[108]  (
    .I(r1do_108_)
  );

zview \I_zview_r1do[107]  (
    .I(r1do_107_)
  );

zview \I_zview_r1do[106]  (
    .I(r1do_106_)
  );

zview \I_zview_r1do[105]  (
    .I(r1do_105_)
  );

zview \I_zview_r1do[104]  (
    .I(r1do_104_)
  );

zview \I_zview_r1do[103]  (
    .I(r1do_103_)
  );

zview \I_zview_r1do[102]  (
    .I(r1do_102_)
  );

zview \I_zview_r1do[101]  (
    .I(r1do_101_)
  );

zview \I_zview_r1do[100]  (
    .I(r1do_100_)
  );

zview \I_zview_r1do[99]  (
    .I(r1do_99_)
  );

zview \I_zview_r1do[98]  (
    .I(r1do_98_)
  );

zview \I_zview_r1do[97]  (
    .I(r1do_97_)
  );

zview \I_zview_r1do[96]  (
    .I(r1do_96_)
  );

zview \I_zview_r1do[95]  (
    .I(r1do_95_)
  );

zview \I_zview_r1do[94]  (
    .I(r1do_94_)
  );

zview \I_zview_r1do[93]  (
    .I(r1do_93_)
  );

zview \I_zview_r1do[92]  (
    .I(r1do_92_)
  );

zview \I_zview_r1do[91]  (
    .I(r1do_91_)
  );

zview \I_zview_r1do[90]  (
    .I(r1do_90_)
  );

zview \I_zview_r1do[89]  (
    .I(r1do_89_)
  );

zview \I_zview_r1do[88]  (
    .I(r1do_88_)
  );

zview \I_zview_r1do[87]  (
    .I(r1do_87_)
  );

zview \I_zview_r1do[86]  (
    .I(r1do_86_)
  );

zview \I_zview_r1do[85]  (
    .I(r1do_85_)
  );

zview \I_zview_r1do[84]  (
    .I(r1do_84_)
  );

zview \I_zview_r1do[83]  (
    .I(r1do_83_)
  );

zview \I_zview_r1do[82]  (
    .I(r1do_82_)
  );

zview \I_zview_r1do[81]  (
    .I(r1do_81_)
  );

zview \I_zview_r1do[80]  (
    .I(r1do_80_)
  );

zview \I_zview_r1do[79]  (
    .I(r1do_79_)
  );

zview \I_zview_r1do[78]  (
    .I(r1do_78_)
  );

zview \I_zview_r1do[77]  (
    .I(r1do_77_)
  );

zview \I_zview_r1do[76]  (
    .I(r1do_76_)
  );

zview \I_zview_r1do[75]  (
    .I(r1do_75_)
  );

zview \I_zview_r1do[74]  (
    .I(r1do_74_)
  );

zview \I_zview_r1do[73]  (
    .I(r1do_73_)
  );

zview \I_zview_r1do[72]  (
    .I(r1do_72_)
  );

zview \I_zview_r1do[71]  (
    .I(r1do_71_)
  );

zview \I_zview_r1do[70]  (
    .I(r1do_70_)
  );

zview \I_zview_r1do[69]  (
    .I(r1do_69_)
  );

zview \I_zview_r1do[68]  (
    .I(r1do_68_)
  );

zview \I_zview_r1do[67]  (
    .I(r1do_67_)
  );

zview \I_zview_r1do[66]  (
    .I(r1do_66_)
  );

zview \I_zview_r1do[65]  (
    .I(r1do_65_)
  );

zview \I_zview_r1do[64]  (
    .I(r1do_64_)
  );

zview \I_zview_r1do[63]  (
    .I(r1do_63_)
  );

zview \I_zview_r1do[62]  (
    .I(r1do_62_)
  );

zview \I_zview_r1do[61]  (
    .I(r1do_61_)
  );

zview \I_zview_r1do[60]  (
    .I(r1do_60_)
  );

zview \I_zview_r1do[59]  (
    .I(r1do_59_)
  );

zview \I_zview_r1do[58]  (
    .I(r1do_58_)
  );

zview \I_zview_r1do[57]  (
    .I(r1do_57_)
  );

zview \I_zview_r1do[56]  (
    .I(r1do_56_)
  );

zview \I_zview_r1do[55]  (
    .I(r1do_55_)
  );

zview \I_zview_r1do[54]  (
    .I(r1do_54_)
  );

zview \I_zview_r1do[53]  (
    .I(r1do_53_)
  );

zview \I_zview_r1do[52]  (
    .I(r1do_52_)
  );

zview \I_zview_r1do[51]  (
    .I(r1do_51_)
  );

zview \I_zview_r1do[50]  (
    .I(r1do_50_)
  );

zview \I_zview_r1do[49]  (
    .I(r1do_49_)
  );

zview \I_zview_r1do[48]  (
    .I(r1do_48_)
  );

zview \I_zview_r1do[47]  (
    .I(r1do_47_)
  );

zview \I_zview_r1do[46]  (
    .I(r1do_46_)
  );

zview \I_zview_r1do[45]  (
    .I(r1do_45_)
  );

zview \I_zview_r1do[44]  (
    .I(r1do_44_)
  );

zview \I_zview_r1do[43]  (
    .I(r1do_43_)
  );

zview \I_zview_r1do[42]  (
    .I(r1do_42_)
  );

zview \I_zview_r1do[41]  (
    .I(r1do_41_)
  );

zview \I_zview_r1do[40]  (
    .I(r1do_40_)
  );

zview \I_zview_r1do[39]  (
    .I(r1do_39_)
  );

zview \I_zview_r1do[38]  (
    .I(r1do_38_)
  );

zview \I_zview_r1do[37]  (
    .I(r1do_37_)
  );

zview \I_zview_r1do[36]  (
    .I(r1do_36_)
  );

zview \I_zview_r1do[35]  (
    .I(r1do_35_)
  );

zview \I_zview_r1do[34]  (
    .I(r1do_34_)
  );

zview \I_zview_r1do[33]  (
    .I(r1do_33_)
  );

zview \I_zview_r1do[32]  (
    .I(r1do_32_)
  );

zview \I_zview_r1do[31]  (
    .I(r1do_31_)
  );

zview \I_zview_r1do[30]  (
    .I(r1do_30_)
  );

zview \I_zview_r1do[29]  (
    .I(r1do_29_)
  );

zview \I_zview_r1do[28]  (
    .I(r1do_28_)
  );

zview \I_zview_r1do[27]  (
    .I(r1do_27_)
  );

zview \I_zview_r1do[26]  (
    .I(r1do_26_)
  );

zview \I_zview_r1do[25]  (
    .I(r1do_25_)
  );

zview \I_zview_r1do[24]  (
    .I(r1do_24_)
  );

zview \I_zview_r1do[23]  (
    .I(r1do_23_)
  );

zview \I_zview_r1do[22]  (
    .I(r1do_22_)
  );

zview \I_zview_r1do[21]  (
    .I(r1do_21_)
  );

zview \I_zview_r1do[20]  (
    .I(r1do_20_)
  );

zview \I_zview_r1do[19]  (
    .I(r1do_19_)
  );

zview \I_zview_r1do[18]  (
    .I(r1do_18_)
  );

zview \I_zview_r1do[17]  (
    .I(r1do_17_)
  );

zview \I_zview_r1do[16]  (
    .I(r1do_16_)
  );

zview \I_zview_r1do[15]  (
    .I(r1do_15_)
  );

zview \I_zview_r1do[14]  (
    .I(r1do_14_)
  );

zview \I_zview_r1do[13]  (
    .I(r1do_13_)
  );

zview \I_zview_r1do[12]  (
    .I(r1do_12_)
  );

zview \I_zview_r1do[11]  (
    .I(r1do_11_)
  );

zview \I_zview_r1do[10]  (
    .I(r1do_10_)
  );

zview \I_zview_r1do[9]  (
    .I(r1do_9_)
  );

zview \I_zview_r1do[8]  (
    .I(r1do_8_)
  );

zview \I_zview_r1do[7]  (
    .I(r1do_7_)
  );

zview \I_zview_r1do[6]  (
    .I(r1do_6_)
  );

zview \I_zview_r1do[5]  (
    .I(r1do_5_)
  );

zview \I_zview_r1do[4]  (
    .I(r1do_4_)
  );

zview \I_zview_r1do[3]  (
    .I(r1do_3_)
  );

zview \I_zview_r1do[2]  (
    .I(r1do_2_)
  );

zview \I_zview_r1do[1]  (
    .I(r1do_1_)
  );

zview \I_zview_r1do[0]  (
    .I(r1do_0_)
  );

endmodule

